** Profile: "SCHEMATIC1-bka"  [ g:\hiast\4th year\second term\����\pspice\trgen-schematic1-bka.sim ] 

** Creating circuit file "trgen-schematic1-bka.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 15m 0 100n SKIPBP 
.OPTIONS ABSTOL= 1.0n
.OPTIONS CHGTOL= 0.01n
.OPTIONS ITL4= 100
.OPTIONS RELTOL= 0.01
.OPTIONS VNTOL= 1.0m
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\trgen-SCHEMATIC1.net" 


.END
