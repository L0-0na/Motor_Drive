** Profile: "SCHEMATIC1-clipper"  [ G:\HIAST\4th year\second term\����\clippers-SCHEMATIC1-clipper.sim ] 

** Creating circuit file "clippers-SCHEMATIC1-clipper.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.4ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\clippers-SCHEMATIC1.net" 


.END
